-- megafunction wizard: %ALTACCUMULATE%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altaccumulate 

-- ============================================================
-- File Name: A.vhd
-- Megafunction Name(s):
-- 			altaccumulate
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.0 Build 184 04/29/2009 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2009 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY A IS
	PORT
	(
		aclr		: IN STD_LOGIC  := '0';
		clken		: IN STD_LOGIC  := '1';
		clock		: IN STD_LOGIC  := '0';
		data		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (4 DOWNTO 0)
	);
END A;


ARCHITECTURE SYN OF a IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (4 DOWNTO 0);



	COMPONENT altaccumulate
	GENERIC (
		lpm_representation		: STRING;
		lpm_type		: STRING;
		width_in		: NATURAL;
		width_out		: NATURAL
	);
	PORT (
			clken	: IN STD_LOGIC ;
			aclr	: IN STD_LOGIC ;
			clock	: IN STD_LOGIC ;
			data	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (4 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(4 DOWNTO 0);

	altaccumulate_component : altaccumulate
	GENERIC MAP (
		lpm_representation => "UNSIGNED",
		lpm_type => "altaccumulate",
		width_in => 4,
		width_out => 5
	)
	PORT MAP (
		clken => clken,
		aclr => aclr,
		clock => clock,
		data => data,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ACLR NUMERIC "1"
-- Retrieval info: PRIVATE: ADD_SUB NUMERIC "0"
-- Retrieval info: PRIVATE: CIN NUMERIC "0"
-- Retrieval info: PRIVATE: CLKEN NUMERIC "1"
-- Retrieval info: PRIVATE: COUT NUMERIC "0"
-- Retrieval info: PRIVATE: EXTRA_LATENCY NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "ACEX1K"
-- Retrieval info: PRIVATE: LATENCY NUMERIC "0"
-- Retrieval info: PRIVATE: LPM_REPRESENTATION NUMERIC "1"
-- Retrieval info: PRIVATE: OVERFLOW NUMERIC "0"
-- Retrieval info: PRIVATE: SLOAD NUMERIC "0"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: WIDTH_IN NUMERIC "4"
-- Retrieval info: PRIVATE: WIDTH_OUT NUMERIC "5"
-- Retrieval info: CONSTANT: LPM_REPRESENTATION STRING "UNSIGNED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altaccumulate"
-- Retrieval info: CONSTANT: WIDTH_IN NUMERIC "4"
-- Retrieval info: CONSTANT: WIDTH_OUT NUMERIC "5"
-- Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT GND aclr
-- Retrieval info: USED_PORT: clken 0 0 0 0 INPUT VCC clken
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT GND clock
-- Retrieval info: USED_PORT: data 0 0 4 0 INPUT NODEFVAL data[3..0]
-- Retrieval info: USED_PORT: result 0 0 5 0 OUTPUT NODEFVAL result[4..0]
-- Retrieval info: CONNECT: @data 0 0 4 0 data 0 0 4 0
-- Retrieval info: CONNECT: result 0 0 5 0 @result 0 0 5 0
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @clken 0 0 0 0 clken 0 0 0 0
-- Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL A.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL A.inc TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL A.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL A.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL A_inst.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL A_waveforms.html TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL A_wave*.jpg FALSE
-- Retrieval info: LIB_FILE: altera_mf
