ComparadorFinal_inst : ComparadorFinal PORT MAP (
		clken	 => clken_sig,
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		AeB	 => AeB_sig,
		AgB	 => AgB_sig,
		AlB	 => AlB_sig
	);
