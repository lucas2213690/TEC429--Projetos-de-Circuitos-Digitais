Comparador21_inst : Comparador21 PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		AeB	 => AeB_sig,
		AgB	 => AgB_sig
	);
