Comparador17_inst : Comparador17 PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		AgeB	 => AgeB_sig
	);
